`timescale 1ns / 1ps

// Inst_Mem��ָ��洢����ֻ����
// - addr Ϊ�ֽڵ�ַ
// - �ڲ����ֶ��룺�� addr[4:2] ѡ�� 8 ��ָ��
module Inst_Mem(
    input [31:0] addr,
    output reg [31:0] inst
);

reg [31:0] inst_mem[0:7];

// initial�������ʼ���̶�ָ������
// Ŀ�ģ���֤ addi/beq/bne/jal/jr/j �Ŀ�������ת
initial begin
    // ����ָ�����У��ȸ�ֵ��beq��bne��jal��jr��j
    inst_mem[0] = 32'h20010005; // addi $1,$0,5 ��$1=5��
    inst_mem[1] = 32'h20020006; // addi $2,$0,6 ��$2=6��ȷ��bne������
    inst_mem[2] = 32'h00010814; // beq $0,$1,4   ��$0��$1������֧��PC+4��0x10��
    inst_mem[3] = 32'h00410815; // bne $2,$1,4   ��$2��$1����֧��0x1C��
    inst_mem[4] = 32'h0c000007; // jal 0x1C      ����ת��д$31=0x14��
    inst_mem[5] = 32'h00000000; // NOP
    inst_mem[6] = 32'h03e00008; // jr $31        ������$31=0x14��
    inst_mem[7] = 32'h08000000; // j 0x0         ���������0x0��
end

// ��϶������� addr[4:2] �����Ӧָ��
always @(*) begin
    case(addr[4:2])
        3'b000: inst = inst_mem[0];
        3'b001: inst = inst_mem[1];
        3'b010: inst = inst_mem[2];
        3'b011: inst = inst_mem[3];
        3'b100: inst = inst_mem[4];
        3'b101: inst = inst_mem[5];
        3'b110: inst = inst_mem[6];
        3'b111: inst = inst_mem[7];
        default: inst = 32'h00000000;
    endcase
end

endmodule