`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Data_Mem�����ݴ洢����RAM ���
// - д��posedge clk ͬ��д��we=1 ʱд��
// - ������϶� always @(*)
// - addr ʹ���ֽڵ�ַ���ڲ�ͨ�� addr[6:2] ӳ��Ϊ word ����
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:53:23 12/02/2025 
// Design Name: 
// Module Name:    Data_Mem 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
// Data_Memģ��������
`timescale 1ns / 1ps

module Data_Mem(
    input clk,          // ʱ��
    input we,           // дʹ�ܣ�����Ч��
    input [31:0] addr,  // 32λ��ַ����
    input [31:0] wr_data, // 32λд����
    output reg [31:0] rd_data // 32λ������
);
    // 1. ģ�鼶�����������ؼ����Ƴ����п飩
    integer i; // ��ʼ���õ���������������ģ�鿪ͷ
    // �������ݴ洢����32��32λ�洢��Ԫ
    reg [31:0] data_mem[0:31]; 

    // 2. ��ʼ�����ݴ洢����ȫ0���޿��ڱ���������
    initial begin
        for(i=0; i<=31; i=i+1) begin
            data_mem[i] = 32'h00000000;
        end
    end

    // 3. д������ʱ���߼���ʱ�������أ�
    //    - we=1 ʱд��
    //    - addr[6:2] ��Ϊ word ����
    always @(posedge clk) begin
        if(we) begin
            case(addr[6:2]) // 5λ��ַƥ��洢��Ԫ
                5'b00000: data_mem[0] = wr_data;
                5'b00001: data_mem[1] = wr_data;
                5'b00010: data_mem[2] = wr_data;
                5'b00011: data_mem[3] = wr_data;
                5'b00100: data_mem[4] = wr_data;
                default: data_mem[0] = wr_data; // Ĭ��д��һ����Ԫ
            endcase
        end
    end

    // 4. ������������߼����޶�̬������
    //    - ֱ�Ӱ� addr[6:2] �����Ӧ data_mem ��
    always @(*) begin
        case(addr[6:2])
            5'b00000: rd_data = data_mem[0];
            5'b00001: rd_data = data_mem[1];
            5'b00010: rd_data = data_mem[2];
            5'b00011: rd_data = data_mem[3];
            5'b00100: rd_data = data_mem[4];
            default: rd_data = 32'h00000000; // �����ַ����0
        endcase
    end

endmodule