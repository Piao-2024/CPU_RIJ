`timescale 1ns / 1ps

// PC�������������Program Counter��
// ���ܣ���ÿ��ʱ�������أ����ݿ����ź� PC_s ѡ����һ��ָ���ַ
//
// PC_s ���루����ע�����Ѷ��壩��
// - 2'b00��˳��ִ�У�PC = PC + 4��
// - 2'b01��jr��PC = R_Data_A��
// - 2'b10����֧��PC = branch_addr��
// - 2'b11����ת��PC = jump_addr��
//
// �ӿ�˵����
// - clk��ʱ�ӣ������ظ��� PC
// - rst_n������Ч�첽��λ��negedge rst_n ������
// - PC_new������˿���д���� PC+4������ǰʵ�ֲ�δʹ�ø����루PC+4��ģ���ڲ����㣩
// - R_Data_A���Ĵ��� rs �Ķ����ݣ����� jr
// - branch_addr����֧Ŀ���ַ��beq/bne �����ⲿ����ã�
// - jump_addr��j/jal Ŀ���ַ�������ⲿƴ��/����ã�
// - PC����ǰ PC���Ĵ�����
// - PC_new_out�������PC+4������ǰʵ��Ϊ�Ĵ��������
module PC(
    input clk,
    input rst_n,
    input [1:0] PC_s,          // PC ѡ���ź�
    input [31:0] R_Data_A,     // jr��PC = rs_data
    input [31:0] branch_addr,  // ��֧Ŀ���ַ
    input [31:0] jump_addr,    // ��תĿ���ַ
    output reg [31:0] PC,      // ��ǰ PC���Ĵ�����
    output [31:0] PC_new_out   // ��� PC+4������߼���ʼ�յ��� PC+4��
);

    // ��������PC_new_out ��Զ��ӳ����ǰ PC + 4��
    // ���� CPU_TOP �ڼ��� branch/jump/jal ��ص�ַʱ��������֡���һ�� PC+4����ʱ���λ��
    assign PC_new_out = PC + 32'h0000_0004;

    always @(posedge clk or negedge rst_n) begin
        if(!rst_n) begin
            // ��λ��PC �� 0 ��ʼȡָ
            PC <= 32'h00000000;
        end else begin
            // ���� PC_s ѡ����һ�� PC ����Դ
            case(PC_s)
                2'b00: PC <= PC + 32'h0000_0004; // ˳��ִ�У�PC = PC + 4
                2'b01: PC <= R_Data_A;    // jr��PC = rs_data
                2'b10: PC <= branch_addr; // ��֧��PC = branch_addr
                2'b11: PC <= jump_addr;   // ��ת��PC = jump_addr
                default: PC <= PC + 32'h0000_0004;
            endcase
        end
    end

endmodule