`timescale 1ns / 1ps

// Controller��������/������
// ���ܣ�����ָ���ֶ� (op/func) ��ȽϽ�� (Zero)��������������ͨ·����Ŀ����ź�
//
// ��Ҫ����ź����壨����㹤������ģ�������ƶϣ���
// - PC_s[1:0]��PC ������Դѡ�񣨼� PC.v��
// - ALU_OP[2:0]��ALU ����ѡ������ 000=add, 001=sub ... ������ ALU ģ��Ϊ׼��
// - imm_s��ALU �ڶ�������ѡ��0=�Ĵ���rt���ݣ�1=��������չֵ��
// - w_r_s[1:0]��д��Ŀ�ļĴ���ѡ��
//   ����00=rd��R�ͣ���01=rt��I�ͣ��� addi����11=$31��jal������������ RegDst/д��ַMUXΪ׼
// - wr_data_s1/wr_data_s0��д������ѡ����λѡ�񣬵ȼ��� wr_data_sel[1:0]��
//   ����jal ��Ҫд PC+4 �� $31����˻�����ĳ�֡�ѡ�� PC+4 ��ͨ����
// - Write_Reg���Ĵ�����дʹ��
// - Mem_Write�����ݴ洢��дʹ�ܣ���ʵ��δʹ��/��δʵ�� sw����˱��� 0��
//
// ˵������ģ���Ǵ�����߼�������仯��������ӳ���������ʱ�ӣ�
module Controller(
    input [5:0] op,
    input [5:0] func,
    input Zero,              // ALU �� Zero ��־�������� beq/bne��
    output reg [1:0] w_r_s,  // д��Ŀ�ļĴ���ѡ��
    output reg imm_s,        // ALU �ڶ�������ѡ�񣨼Ĵ���/��������
    output reg wr_data_s1,   // д������ѡ�� bit1
    output reg wr_data_s0,   // д������ѡ�� bit0
    output reg [2:0] ALU_OP, // ALU ���������
    output reg Write_Reg,    // �Ĵ���дʹ��
    output reg Mem_Write,    // ���ݴ洢��дʹ��
    output reg [1:0] PC_s    // PC ������Դѡ��
);

always @(*) begin
    // =========================================================
    // 1) Ĭ��ֵ����ȫ̬��
    // δʶ��ָ��ʱ��
    // - ��д�Ĵ���
    // - ��д�ڴ�
    // - PC Ĭ��˳��ִ�� +4
    // =========================================================
    w_r_s      = 2'b00;
    imm_s      = 1'b0;
    wr_data_s1 = 1'b0;
    wr_data_s0 = 1'b0;
    ALU_OP     = 3'b000;
    Write_Reg  = 1'b0;
    Mem_Write  = 1'b0;
    PC_s       = 2'b00;

    // =========================================================
    // 2) �����룺�� opcode ����ָ������
    // =========================================================
    case(op)
        // -----------------------------------------------------
        // R �ͣ�����ֻʵ�� jr��func=001000��
        // -----------------------------------------------------
        6'b000000: begin    
            case(func)
                6'b001000: begin // jr rs
                    // jr ��д�Ĵ�����ֻ�ı� PC
                    PC_s      = 2'b01; // PC = R_Data_A
                    Write_Reg = 1'b0;
                end
                default: begin
                    // ���� R ��δʵ�֣�����Ĭ�ϰ�ȫ̬
                end
            endcase
        end

        // -----------------------------------------------------
        // beq���� rs == rt ���֧
        // ����ʵ�֣�ALU �� rs - rt�������Ϊ 0 �� Zero=1
        // -----------------------------------------------------
        6'b000100: begin // beq rs,rt,label
            imm_s  = 1'b0;     // ALU �ڶ��������üĴ���rt�����ڱȽ� rs �� rt��
            ALU_OP = 3'b001;   // sub������ 001 ��ʾ������
            PC_s   = Zero ? 2'b10 : 2'b00; // Zero=1 ��ѡ�� branch_addr������ PC+4
            Write_Reg = 1'b0;  // beq ��д�Ĵ���
        end

        // -----------------------------------------------------
        // bne���� rs != rt ���֧
        // -----------------------------------------------------
        6'b000101: begin // bne rs,rt,label
            imm_s  = 1'b0;
            ALU_OP = 3'b001;   // sub
            PC_s   = (!Zero) ? 2'b10 : 2'b00; // Zero=0 �ŷ�֧
            Write_Reg = 1'b0;
        end

        // -----------------------------------------------------
        // j����������ת
        // -----------------------------------------------------
        6'b000010: begin // j label
            PC_s      = 2'b11; // PC = jump_addr
            Write_Reg = 1'b0;
        end

        // -----------------------------------------------------
        // jal����ת������
        // - PC ��ת�� jump_addr
        // - ͬʱ�ѡ����ص�ַ PC+4��д�� $31
        // -----------------------------------------------------
        6'b000011: begin // jal label
            PC_s      = 2'b11; // ��ת
            w_r_s     = 2'b11; // Ŀ�ļĴ���ѡ�� $31
            wr_data_s1= 1'b1;  // д������ѡ��PC+4���������ȡ������д��MUX��
            wr_data_s0= 1'b0;  // ����/������ 2'b10 �� 2'b??����������ͨ·���壩
            Write_Reg = 1'b1;  // ����д�� $31
        end

        // -----------------------------------------------------
        // addi��rt = rs + signext(imm)
        // ���ڳ�ʼ���Ĵ���ֵ�����ں�����֧�Ƚ�
        // -----------------------------------------------------
        6'b001000: begin // addi rt,rs,offset
            imm_s     = 1'b1;    // ALU �ڶ���������������
            ALU_OP    = 3'b000;  // add������ 000 ��ʾ�ӷ���
            w_r_s     = 2'b01;   // Ŀ�ļĴ���ѡ�� rt
            Write_Reg = 1'b1;    // д�ؽ�����Ĵ���
            PC_s      = 2'b00;   // ���� +4
        end

        default: begin
            // δʵ��ָ�����Ĭ�ϰ�ȫ̬
        end
    endcase
end

endmodule