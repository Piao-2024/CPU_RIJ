`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Data_Mem�����ݴ洢������ RAM��
//
// ���ԣ�
// - д��ͬ��д��posedge clk����we=1 ʱд��
// - ������϶���always @(*)������ַ�仯������ӳ�� rd_data
// - addr���ֽڵ�ַ��byte address��
//   �ڲ��� addr[6:2] ��Ϊ word ������
//   - [1:0] �����ԣ��ȼ��� word ���룩
//   - [6:2] �ɱ�ʾ 0~31��32 �� word��
//
// ע�⣺��ǰ case ֻʵ���� 0~4 �ĵ�ַӳ�䣺
// - ����������ַĬ����� 0
// - д��������ַĬ��д�� data_mem[0]
// ������ƿ��õ�ַ��Χ�����ڡ�ʵ��򻯰汾������Ϊ
//////////////////////////////////////////////////////////////////////////////////

module Data_Mem(
    input clk,             // ʱ�ӣ�д����������Ч
    input we,              // дʹ�ܣ�����Ч��
    input [31:0] addr,     // �ֽڵ�ַ
    input [31:0] wr_data,  // д������
    output reg [31:0] rd_data // �������ݣ��������Ĵ�����
);

    // ��ʼ��ѭ���ñ���������������ģ��������Verilog �﷨Ҫ��
    integer i;

    // 32 x 32-bit �洢���У�word addressed��
    reg [31:0] data_mem[0:31];

    // ��ʼ��������ʱ�� RAM ���㣨�ۺϵ� FPGA ʱ�����ƶϳɳ�ʼ���򱻺��ԣ��ӹ�����������
    initial begin
        for(i=0; i<=31; i=i+1) begin
            data_mem[i] = 32'h00000000;
        end
    end

    // =========================================================
    // д������ͬ��д��posedge clk��
    // =========================================================
    always @(posedge clk) begin
        if(we) begin
            // �� addr[6:2] ��Ϊ word �������ȼ� addr/4��
            case(addr[6:2])
                5'b00000: data_mem[0] <= wr_data;
                5'b00001: data_mem[1] <= wr_data;
                5'b00010: data_mem[2] <= wr_data;
                5'b00011: data_mem[3] <= wr_data;
                5'b00100: data_mem[4] <= wr_data;

                // ������ַ����ǰʵ��д�� 0 �ŵ�Ԫ����/ռλ��Ϊ��
                default:  data_mem[0] <= wr_data;
            endcase
        end
    end

    // =========================================================
    // ����������϶�����ַ�仯�������������
    // =========================================================
    always @(*) begin
        case(addr[6:2])
            5'b00000: rd_data = data_mem[0];
            5'b00001: rd_data = data_mem[1];
            5'b00010: rd_data = data_mem[2];
            5'b00011: rd_data = data_mem[3];
            5'b00100: rd_data = data_mem[4];

            // ������ַ������ 0����/ռλ��Ϊ��
            default:  rd_data = 32'h00000000;
        endcase
    end

endmodule