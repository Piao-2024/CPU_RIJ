`timescale 1ns / 1ps

// Reg_File���Ĵ����ѣ�32��32��
// - д��posedge clk �� Write_Reg=1 ʱд��
// - ������϶���always @(*)��
// - Լ����$0 ��Ϊ 0������ַΪ 0 ʱǿ����� 0��
module Reg_File(
    input clk,
    input rst_n,
    input Write_Reg,
    input [4:0] rs_addr,
    input [4:0] rt_addr,
    input [4:0] rd_addr,
    input [1:0] w_r_s,      // д��ַѡ�񣨽̲�w_r_s��
    input [31:0] wr_data,
    output reg [31:0] rs_data,
    output reg [31:0] rt_data,
    output [31:0] R1_out,   // ����$1�������ȡ
    output [31:0] R31_out   // ����$31�������ȡ
);

reg [31:0] regs[0:31]; // �ڲ��Ĵ������飨reg���ͣ�
integer i;

// ��λ��д�Ĵ���
// - rst_n=0������ȫ���Ĵ���
// - Write_Reg=1������ w_r_s ѡ��д rd/rt/$31
always @(posedge clk or negedge rst_n) begin
    if(!rst_n) begin
        for(i=0; i<=31; i=i+1) regs[i] <= 32'h00000000;
    end else if(Write_Reg) begin
        case(w_r_s)
            2'b11: regs[31] <= wr_data; // jalд$31
            2'b01: regs[rt_addr] <= wr_data;
            2'b00: regs[rd_addr] <= wr_data;
            default: ;
        endcase
    end
end

// ���Ĵ���
// - ���� $0����ַ 0����������� 0
always @(*) begin
    rs_data = (rs_addr == 5'd0) ? 32'h00000000 : regs[rs_addr];
    rt_data = (rt_addr == 5'd0) ? 32'h00000000 : regs[rt_addr];
end

// ����ָ���Ĵ���ֵ����wire��ת������ֱ��assign reg���飩
wire [31:0] R1;
wire [31:0] R31;
assign R1 = regs[1];       // reg����ֵ����wire���Ϸ���
assign R31 = regs[31];
assign R1_out = R1;        // �˿ڵ���wireֵ
assign R31_out = R31;

endmodule