`timescale 1ns / 1ps

// CPU_TB������ƽ̨
// - ����ʱ�� clk��20ns ���ڣ�
// - ������λ rst_n������Ч��
// - ��ӡ CPU_TOP �����Ĺؼ��ź�
module CPU_TB;

reg clk;
reg rst_n;
wire [31:0] PC_out;
wire [31:0] Inst_out;
wire [31:0] ALU_Out_out;
wire Zero_out;
wire [31:0] R1_out;
wire [31:0] R31_out;

// ��������ģ��
CPU_TOP cpu(
    .clk(clk),
    .rst_n(rst_n),
    .PC_out(PC_out),
    .Inst_out(Inst_out),
    .ALU_Out_out(ALU_Out_out),
    .Zero_out(Zero_out),
    .R1_out(R1_out),
    .R31_out(R31_out)
);

// ʱ�����ɣ�20ns���ڣ�
initial begin
    clk = 0;
    forever #10 clk = ~clk;
end

// ��λ�ź�
initial begin
    rst_n = 0;
    #15 rst_n = 1;
end

// ��ӡ���Խ��
// $display����ӡһ��
// $monitor���źű仯����ӡ
initial begin
    $display("------------------------ʵ��ָ�����------------------------");
    $monitor("Time=%0d | PC=%h | Inst=%h | ALU_Out=%h | Zero=%b | R1=%h | R31=%h",
        $time, PC_out, Inst_out, ALU_Out_out, Zero_out, R1_out, R31_out);
    #1000 $stop;
end

endmodule