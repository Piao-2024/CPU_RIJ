`timescale 1ns / 1ps

// PC�����������
// - PC_s=00��˳��ִ�У�PC+4��
// - PC_s=01��jr��PC=rs_data��
// - PC_s=10����֧��PC=branch_addr��
// - PC_s=11����ת��PC=jump_addr��
module PC(
    input clk,
    input rst_n,
    input [1:0] PC_s,       // �̲ı�14.26��PC_s
    input [31:0] PC_new,    // PC+4
    input [31:0] R_Data_A,  // rs_data��jrָ�
    input [31:0] branch_addr, // ��֧��ַ��beq/bne��
    input [31:0] jump_addr,  // J����ת��ַ��j/jal��
    output reg [31:0] PC,   // ��ǰPC
    output reg [31:0] PC_new_out // PC+4�������Ϊreg��
);

// ʱ���߼�����ʱ���ظ��� PC������� PC+4
// ��λ��rst_n=0 ʱ PC �� 0
always @(posedge clk or negedge rst_n) begin
    if(!rst_n) begin
        PC <= 32'h00000000;
        PC_new_out <= 32'h00000004;
    end else begin
        PC_new_out <= PC + 32'h00000004; // ʱ���ظ���PC+4
        case(PC_s)
            2'b00: PC <= PC_new_out;        // ����+4
            2'b01: PC <= R_Data_A;          // jrָ�rs_data��
            2'b10: PC <= branch_addr;       // beq/bne��֧
            2'b11: PC <= jump_addr;         // j/jal��ת
        endcase
    end
end

endmodule