`timescale 1ns / 1ps

// Controller��������/������
// - ���룺op/func��ָ���ֶΣ���Zero��ALU �ȽϽ����
// - �����PC_s / ALU_OP / imm_s / Write_Reg / w_r_s / wr_data_s* / Mem_Write
module Controller(
    input [5:0] op,
    input [5:0] func,
    input Zero,             // ALU���־��beq/bne�жϣ�
    output reg [1:0] w_r_s, // д��ַѡ��
    output reg imm_s,       // ALUԴѡ��
    output reg wr_data_s1,  // д����ѡ��λ1
    output reg wr_data_s0,  // д����ѡ��λ0
    output reg [2:0] ALU_OP,// ALU������
    output reg Write_Reg,   // �Ĵ���дʹ��
    output reg Mem_Write,   // �洢��дʹ�ܣ�ʵ��δҪ����0��
    output reg [1:0] PC_s   // PCѡ���ź�
);

always @(*) begin
    // Ĭ��ֵ��ʼ����δʶ��ָ��ʱ�ġ���ȫ̬����
    // - PC_s=00��˳��ִ�У�PC+4��
    // - Write_Reg/Mem_Write=0����д�Ĵ���/��д�ڴ�
    w_r_s = 2'b00;
    imm_s = 1'b0;
    wr_data_s1 = 1'b0;
    wr_data_s0 = 1'b0;
    ALU_OP = 3'b000;
    Write_Reg = 1'b0;
    Mem_Write = 1'b0;
    PC_s = 2'b00; // Ĭ��PC+4

    // op ����
    case(op)
        6'b000000: begin // R��ָ���ʵ��jr��
            // func ��һ������
            case(func)
                6'b001000: begin // jr rs
                    PC_s = 2'b01; // ѡrs_data��ΪPC
                    Write_Reg = 1'b0;
                end
                default: ;
            endcase
        end
        6'b000100: begin // beq rs,rt,label
            imm_s = 1'b0;
            ALU_OP = 3'b001; // ALU������
            PC_s = Zero ? 2'b10 : 2'b00; // Zero=1���֧
            Write_Reg = 1'b0;
        end
        6'b000101: begin // bne rs,rt,label
            imm_s = 1'b0;
            ALU_OP = 3'b001; // ALU������
            PC_s = !Zero ? 2'b10 : 2'b00; // Zero=0���֧
            Write_Reg = 1'b0;
        end
        6'b000010: begin // j label
            PC_s = 2'b11; // ѡJ����ת��ַ
            Write_Reg = 1'b0;
        end
        6'b000011: begin // jal label
            PC_s = 2'b11; // ѡJ����ת��ַ
            w_r_s = 2'b11; // д$31��ra��
            wr_data_s1 = 1'b1; // д����ΪPC+4
            Write_Reg = 1'b1; // д��$31
        end
        // addi�����ڳ�ʼ���Ĵ���ֵ�����ڷ�֧�Ƚ�
        6'b001000: begin // addi rt,rs,offset
            imm_s = 1'b1;    // ALUԴѡ������
            ALU_OP = 3'b000; // ALU���ӷ�
            w_r_s = 2'b01;   // д��ַѡrt
            Write_Reg = 1'b1;// ����д�Ĵ���
            PC_s = 2'b00;    // PC����+4
        end
        default: ;
    endcase
end

endmodule