`timescale 1ns / 1ps

// ALU????????????
// - ? ALU_OP ??? a?b ???
// - Zero = (ALU_Out == 0)??? beq/bne ???????
module ALU(
    input [31:0] a,
    input [31:0] b,
    input [2:0] ALU_OP,
    output reg [31:0] ALU_Out,
    output reg Zero
);

// ???????????????
always @(*) begin
    // ALU_OP=000????addi?
    // ALU_OP=001????beq/bne ?????????
    // ????? 0
    case(ALU_OP)
        3'b000: ALU_Out = a + b; // �ӷ���addi��
        3'b001: ALU_Out = a - b; // ������beq/bne��
        default: ALU_Out = 32'h00000000;
    endcase

    // Zero ???????? 0
    Zero = (ALU_Out == 32'h00000000) ? 1'b1 : 1'b0;
end

endmodule