`timescale 1ns / 1ps

// CPU_TOP������ģ�飨�������� CPU ����ͨ·��
// ��Ҫ���ӹ�ϵ��
//   PC -> Inst_Mem -> (�ֶβ��) -> Controller/Reg_File/Imm_Ext -> ALU
//   Controller ���������źţ�PC_s/ALU_OP/imm_s/Write_Reg/w_r_s/wr_data_s*
//   Data_Mem ��ʵ���������ߣ�wr_data_s0 ��ѡ��������ݣ����ں�����չ lw��
module CPU_TOP(
    input clk,
    input rst_n,
    // ��TB��ӡ���ź�
    output [31:0] PC_out,
    output [31:0] Inst_out,
    output [31:0] ALU_Out_out,
    output Zero_out,
    output [31:0] R1_out,
    output [31:0] R31_out // $31��ra��������jalָ��
);

// -----------------------------
// �ڲ��źţ�PC/ָ��/�Ĵ���/����/��ַ��
// -----------------------------
// �ڲ��źŶ��壨����Data_Mem����źţ�
wire [31:0] PC;
wire [31:0] PC_new; // PC+4
wire [31:0] Inst;
wire [5:0] op;
wire [5:0] func;
wire [4:0] rs_addr;
wire [4:0] rt_addr;
wire [4:0] rd_addr;
wire [4:0] shamt;
wire [15:0] imm_offset;
wire [25:0] j_addr;
wire [31:0] imm_ext; // ������չ���������
wire [31:0] rs_data;
wire [31:0] rt_data;
wire [31:0] wr_data;
wire [31:0] ALU_Out;
wire Zero;
wire [1:0] PC_s; // PCѡ���ź�
wire [1:0] w_r_s; // д��ַѡ��
wire imm_s;      // ALUԴѡ��
wire wr_data_s1;  // д����ѡ��λ1
wire wr_data_s0;  // д����ѡ��λ0������������ѡ��Data_Mem�����ݣ�
wire [2:0] ALU_OP;
wire Write_Reg;
wire Mem_Write;
wire [31:0] branch_addr; // ��֧��ַ��PC+4 + offset*4��
wire [31:0] jump_addr;   // J����ת��ַ��PC[31:28]+address+2'b00��
wire [31:0] jal_addr;    // jalָ��д�ص�$raֵ��PC+4��
// Data_Mem�����ź�
wire [31:0] data_mem_rd_data; // Data_Mem������
wire [31:0] data_mem_wr_data; // Data_Memд���ݣ�����rt_data��

// -----------------------------
// ��ģ��ʵ������PC / Inst_Mem / Controller / Reg_File / Imm_Ext / ALU / Data_Mem
// -----------------------------

// 1. PCģ��
PC pc_module(
    .clk(clk),
    .rst_n(rst_n),
    .PC_s(PC_s),
    .R_Data_A(rs_data),
    .branch_addr(branch_addr),
    .jump_addr(jump_addr),
    .PC(PC),
    .PC_new_out(PC_new)
);

// ָ��洢����addr=PC -> inst=Inst
// 2. ָ��洢����Inst_Mem��
Inst_Mem inst_mem(
    .addr(PC),
    .inst(Inst)
);

// 3. �����������̲ı�14.26���ɿ����źţ�
Controller ctrl(
    .op(op),
    .func(func),
    .Zero(Zero),
    .w_r_s(w_r_s),
    .imm_s(imm_s),
    .wr_data_s1(wr_data_s1),
    .wr_data_s0(wr_data_s0), // ���ӿ�������wr_data_s0
    .ALU_OP(ALU_OP),
    .Write_Reg(Write_Reg),
    .Mem_Write(Mem_Write),
    .PC_s(PC_s)
);

// �Ĵ����ѣ����� rs_data/rt_data��д���� Write_Reg + w_r_s ����
// 4. �Ĵ����ѣ�֧��$31д�أ�
Reg_File reg_file(
    .clk(clk),
    .rst_n(rst_n),
    .Write_Reg(Write_Reg),
    .rs_addr(rs_addr),
    .rt_addr(rt_addr),
    .rd_addr(rd_addr),
    .w_r_s(w_r_s),
    .wr_data(wr_data),
    .rs_data(rs_data),
    .rt_data(rt_data),
    .R1_out(R1_out),
    .R31_out(R31_out)
);

// ��������չ��Inst[15:0] -> imm_ext��������չ��
// 5. ������������չ
Imm_Ext imm_ext_module(
    .imm(imm_offset),
    .imm_ext(imm_ext)
);

// 6. ALU��ʵ������/�߼�/��λ���㣩
ALU alu_module(
    .a(rs_data),
    .b(imm_s ? imm_ext : rt_data),
    .ALU_OP(ALU_OP),
    .ALU_Out(ALU_Out),
    .Zero(Zero)
);

// ���ݴ洢����addr=ALU_Out��д����=rt_data��������=rd_data���� lw Ԥ����
// 7. ���ݴ洢����Data_Mem��������
Data_Mem data_mem_module(
    .clk(clk),
    .we(Mem_Write),       // дʹ�ܣ��ӿ�������Mem_Write
    .addr(ALU_Out),       // ��ַ��ALU��������lw/sw�ĵ�ַ��
    .wr_data(rt_data),    // д���ݣ��Ĵ����ѵ�rt_data��swָ��Դ���ݣ�
    .rd_data(data_mem_rd_data) // �����ݣ������д��ѡ��
);

// -----------------------------
// ����߼�����֧/��ת��ַ���㡢д������ѡ���ֶβ��
// -----------------------------

// 8. ��ַ���㣨��֧/��ת��
assign branch_addr = PC_new + (imm_ext << 2); // PC+4 + offset*4
assign jump_addr = {PC_new[31:28], j_addr, 2'b00}; // J�͵�ַƴ��
assign jal_addr = PC_new; // jalָ��д��$31�ĵ�ַ��PC+4��

// д������ѡ��
//   wr_data_s1=1 -> jal_addr(PC+4)
//   wr_data_s0=1 -> data_mem_rd_data��Ԥ���� lw��
//   ����         -> ALU_Out������ addi��
// 9. д����ѡ������Data_Mem�����ݵ�ѡ��
assign wr_data = wr_data_s1 ? jal_addr : (wr_data_s0 ? data_mem_rd_data : ALU_Out);

// ָ���ֶ���ȡ
assign op = Inst[31:26];
assign func = Inst[5:0];
assign rs_addr = Inst[25:21];
assign rt_addr = Inst[20:16];
assign rd_addr = Inst[15:11];
assign shamt = Inst[10:6];
assign imm_offset = Inst[15:0];
assign j_addr = Inst[25:0];

// ����˿ڣ���TB��ӡ��
assign PC_out = PC;
assign Inst_out = Inst;
assign ALU_Out_out = ALU_Out;
assign Zero_out = Zero;

endmodule